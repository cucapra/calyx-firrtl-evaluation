module main(
  input         go,
  input         clk,
  input         reset,
  output        done,
  output [3:0]  A_int_addr0,
  output [3:0]  A_int_addr1,
  output        A_int_write_en,
  output [31:0] A_int_write_data,
  output        A_int_read_en,
  input  [31:0] A_int_read_data,
  input         A_int_write_done,
  input         A_int_read_done,
  output [3:0]  B_int_addr0,
  output [3:0]  B_int_addr1,
  output        B_int_write_en,
  output [31:0] B_int_write_data,
  output        B_int_read_en,
  input  [31:0] B_int_read_data,
  input         B_int_write_done,
  input         B_int_read_done,
  output [3:0]  C_int_addr0,
  output [3:0]  C_int_addr1,
  output        C_int_write_en,
  output [31:0] C_int_write_data,
  output        C_int_read_en,
  input  [31:0] C_int_read_data,
  input         C_int_write_done,
  input         C_int_read_done,
  output        alpha_int_addr0,
  output        alpha_int_write_en,
  output [31:0] alpha_int_write_data,
  output        alpha_int_read_en,
  input  [31:0] alpha_int_read_data,
  input         alpha_int_write_done,
  input         alpha_int_read_done,
  output        beta_int_addr0,
  output        beta_int_write_en,
  output [31:0] beta_int_write_data,
  output        beta_int_read_en,
  input  [31:0] beta_int_read_data,
  input         beta_int_write_done,
  input         beta_int_read_done
);
  wire [31:0] A_int_read0_0_in;
  wire  A_int_read0_0_write_en;
  wire  A_int_read0_0_clk;
  wire  A_int_read0_0_reset;
  wire [31:0] A_int_read0_0_out;
  wire  A_int_read0_0_done;
  wire [31:0] B_int_read0_0_in;
  wire  B_int_read0_0_write_en;
  wire  B_int_read0_0_clk;
  wire  B_int_read0_0_reset;
  wire [31:0] B_int_read0_0_out;
  wire  B_int_read0_0_done;
  wire [31:0] C_i_j_0_in;
  wire  C_i_j_0_write_en;
  wire  C_i_j_0_clk;
  wire  C_i_j_0_reset;
  wire [31:0] C_i_j_0_out;
  wire  C_i_j_0_done;
  wire [3:0] add2_left;
  wire [3:0] add2_right;
  wire [3:0] add2_out;
  wire [31:0] add3_left;
  wire [31:0] add3_right;
  wire [31:0] add3_out;
  wire [31:0] add4_left;
  wire [31:0] add4_right;
  wire [31:0] add4_out;
  wire [31:0] alpha_int_read0_0_in;
  wire  alpha_int_read0_0_write_en;
  wire  alpha_int_read0_0_clk;
  wire  alpha_int_read0_0_reset;
  wire [31:0] alpha_int_read0_0_out;
  wire  alpha_int_read0_0_done;
  wire [31:0] beta_int_read0_0_in;
  wire  beta_int_read0_0_write_en;
  wire  beta_int_read0_0_clk;
  wire  beta_int_read0_0_reset;
  wire [31:0] beta_int_read0_0_out;
  wire  beta_int_read0_0_done;
  wire [31:0] const0_out;
  wire [3:0] const1_out;
  wire  const10_out;
  wire [3:0] const11_out;
  wire [3:0] const2_out;
  wire [3:0] const4_out;
  wire  const9_out;
  wire [3:0] i0_in;
  wire  i0_write_en;
  wire  i0_clk;
  wire  i0_reset;
  wire [3:0] i0_out;
  wire  i0_done;
  wire [3:0] j0_in;
  wire  j0_write_en;
  wire  j0_clk;
  wire  j0_reset;
  wire [3:0] j0_out;
  wire  j0_done;
  wire [3:0] k_0_in;
  wire  k_0_write_en;
  wire  k_0_clk;
  wire  k_0_reset;
  wire [3:0] k_0_out;
  wire  k_0_done;
  wire [3:0] le0_left;
  wire [3:0] le0_right;
  wire  le0_out;
  wire [3:0] lt0_left;
  wire [3:0] lt0_right;
  wire  lt0_out;
  wire  mult_pipe0_clk;
  wire  mult_pipe0_reset;
  wire  mult_pipe0_go;
  wire [31:0] mult_pipe0_left;
  wire [31:0] mult_pipe0_right;
  wire [31:0] mult_pipe0_out;
  wire  mult_pipe0_done;
  wire [31:0] temp2_0_in;
  wire  temp2_0_write_en;
  wire  temp2_0_clk;
  wire  temp2_0_reset;
  wire [31:0] temp2_0_out;
  wire  temp2_0_done;
  wire  comb_reg_in;
  wire  comb_reg_write_en;
  wire  comb_reg_clk;
  wire  comb_reg_reset;
  wire  comb_reg_out;
  wire  comb_reg_done;
  wire  comb_reg0_in;
  wire  comb_reg0_write_en;
  wire  comb_reg0_clk;
  wire  comb_reg0_reset;
  wire  comb_reg0_out;
  wire  comb_reg0_done;
  wire  comb_reg1_in;
  wire  comb_reg1_write_en;
  wire  comb_reg1_clk;
  wire  comb_reg1_reset;
  wire  comb_reg1_out;
  wire  comb_reg1_done;
  wire [4:0] fsm_in;
  wire  fsm_write_en;
  wire  fsm_clk;
  wire  fsm_reset;
  wire [4:0] fsm_out;
  wire  fsm_done;
  wire  ud_out;
  wire [4:0] adder_left;
  wire [4:0] adder_right;
  wire [4:0] adder_out;
  wire  ud0_out;
  wire [4:0] adder0_left;
  wire [4:0] adder0_right;
  wire [4:0] adder0_out;
  wire  ud1_out;
  wire [4:0] adder1_left;
  wire [4:0] adder1_right;
  wire [4:0] adder1_out;
  wire  ud2_out;
  wire [4:0] adder2_left;
  wire [4:0] adder2_right;
  wire [4:0] adder2_out;
  wire  ud3_out;
  wire [4:0] adder3_left;
  wire [4:0] adder3_right;
  wire [4:0] adder3_out;
  wire  ud4_out;
  wire [4:0] adder4_left;
  wire [4:0] adder4_right;
  wire [4:0] adder4_out;
  wire  ud5_out;
  wire [4:0] adder5_left;
  wire [4:0] adder5_right;
  wire [4:0] adder5_out;
  wire  ud6_out;
  wire [4:0] adder6_left;
  wire [4:0] adder6_right;
  wire [4:0] adder6_out;
  wire  signal_reg_in;
  wire  signal_reg_write_en;
  wire  signal_reg_clk;
  wire  signal_reg_reset;
  wire  signal_reg_out;
  wire  signal_reg_done;
  wire [1:0] fsm0_in;
  wire  fsm0_write_en;
  wire  fsm0_clk;
  wire  fsm0_reset;
  wire [1:0] fsm0_out;
  wire  fsm0_done;
  wire  pd_in;
  wire  pd_write_en;
  wire  pd_clk;
  wire  pd_reset;
  wire  pd_out;
  wire  pd_done;
  wire [1:0] fsm1_in;
  wire  fsm1_write_en;
  wire  fsm1_clk;
  wire  fsm1_reset;
  wire [1:0] fsm1_out;
  wire  fsm1_done;
  wire  pd0_in;
  wire  pd0_write_en;
  wire  pd0_clk;
  wire  pd0_reset;
  wire  pd0_out;
  wire  pd0_done;
  wire [1:0] fsm2_in;
  wire  fsm2_write_en;
  wire  fsm2_clk;
  wire  fsm2_reset;
  wire [1:0] fsm2_out;
  wire  fsm2_done;
  wire  pd1_in;
  wire  pd1_write_en;
  wire  pd1_clk;
  wire  pd1_reset;
  wire  pd1_out;
  wire  pd1_done;
  wire [1:0] fsm3_in;
  wire  fsm3_write_en;
  wire  fsm3_clk;
  wire  fsm3_reset;
  wire [1:0] fsm3_out;
  wire  fsm3_done;
  wire  pd2_in;
  wire  pd2_write_en;
  wire  pd2_clk;
  wire  pd2_reset;
  wire  pd2_out;
  wire  pd2_done;
  wire [1:0] fsm4_in;
  wire  fsm4_write_en;
  wire  fsm4_clk;
  wire  fsm4_reset;
  wire [1:0] fsm4_out;
  wire  fsm4_done;
  wire  pd3_in;
  wire  pd3_write_en;
  wire  pd3_clk;
  wire  pd3_reset;
  wire  pd3_out;
  wire  pd3_done;
  wire [1:0] fsm5_in;
  wire  fsm5_write_en;
  wire  fsm5_clk;
  wire  fsm5_reset;
  wire [1:0] fsm5_out;
  wire  fsm5_done;
  wire  pd4_in;
  wire  pd4_write_en;
  wire  pd4_clk;
  wire  pd4_reset;
  wire  pd4_out;
  wire  pd4_done;
  wire [1:0] fsm6_in;
  wire  fsm6_write_en;
  wire  fsm6_clk;
  wire  fsm6_reset;
  wire [1:0] fsm6_out;
  wire  fsm6_done;
  wire  pd5_in;
  wire  pd5_write_en;
  wire  pd5_clk;
  wire  pd5_reset;
  wire  pd5_out;
  wire  pd5_done;
  wire [1:0] fsm7_in;
  wire  fsm7_write_en;
  wire  fsm7_clk;
  wire  fsm7_reset;
  wire [1:0] fsm7_out;
  wire  fsm7_done;
  wire  pd6_in;
  wire  pd6_write_en;
  wire  pd6_clk;
  wire  pd6_reset;
  wire  pd6_out;
  wire  pd6_done;
  wire [1:0] fsm8_in;
  wire  fsm8_write_en;
  wire  fsm8_clk;
  wire  fsm8_reset;
  wire [1:0] fsm8_out;
  wire  fsm8_done;
  wire  pd7_in;
  wire  pd7_write_en;
  wire  pd7_clk;
  wire  pd7_reset;
  wire  pd7_out;
  wire  pd7_done;
  wire [4:0] fsm9_in;
  wire  fsm9_write_en;
  wire  fsm9_clk;
  wire  fsm9_reset;
  wire [4:0] fsm9_out;
  wire  fsm9_done;
  wire  beg_spl_let10_go_in;
  wire  beg_spl_let10_go_out;
  wire  beg_spl_let10_done_in;
  wire  beg_spl_let10_done_out;
  wire  beg_spl_let11_go_in;
  wire  beg_spl_let11_go_out;
  wire  beg_spl_let11_done_in;
  wire  beg_spl_let11_done_out;
  wire  beg_spl_let13_go_in;
  wire  beg_spl_let13_go_out;
  wire  beg_spl_let13_done_in;
  wire  beg_spl_let13_done_out;
  wire  beg_spl_let14_go_in;
  wire  beg_spl_let14_go_out;
  wire  beg_spl_let14_done_in;
  wire  beg_spl_let14_done_out;
  wire  beg_spl_let15_go_in;
  wire  beg_spl_let15_go_out;
  wire  beg_spl_let15_done_in;
  wire  beg_spl_let15_done_out;
  wire  beg_spl_let16_go_in;
  wire  beg_spl_let16_go_out;
  wire  beg_spl_let16_done_in;
  wire  beg_spl_let16_done_out;
  wire  beg_spl_let17_go_in;
  wire  beg_spl_let17_go_out;
  wire  beg_spl_let17_done_in;
  wire  beg_spl_let17_done_out;
  wire  beg_spl_let4_go_in;
  wire  beg_spl_let4_go_out;
  wire  beg_spl_let4_done_in;
  wire  beg_spl_let4_done_out;
  wire  beg_spl_let5_go_in;
  wire  beg_spl_let5_go_out;
  wire  beg_spl_let5_done_in;
  wire  beg_spl_let5_done_out;
  wire  beg_spl_let6_go_in;
  wire  beg_spl_let6_go_out;
  wire  beg_spl_let6_done_in;
  wire  beg_spl_let6_done_out;
  wire  beg_spl_let7_go_in;
  wire  beg_spl_let7_go_out;
  wire  beg_spl_let7_done_in;
  wire  beg_spl_let7_done_out;
  wire  invoke2_go_in;
  wire  invoke2_go_out;
  wire  invoke2_done_in;
  wire  invoke2_done_out;
  wire  invoke5_go_in;
  wire  invoke5_go_out;
  wire  invoke5_done_in;
  wire  invoke5_done_out;
  wire  invoke6_go_in;
  wire  invoke6_go_out;
  wire  invoke6_done_in;
  wire  invoke6_done_out;
  wire  invoke7_go_in;
  wire  invoke7_go_out;
  wire  invoke7_done_in;
  wire  invoke7_done_out;
  wire  invoke8_go_in;
  wire  invoke8_go_out;
  wire  invoke8_done_in;
  wire  invoke8_done_out;
  wire  invoke13_go_in;
  wire  invoke13_go_out;
  wire  invoke13_done_in;
  wire  invoke13_done_out;
  wire  invoke14_go_in;
  wire  invoke14_go_out;
  wire  invoke14_done_in;
  wire  invoke14_done_out;
  wire  invoke19_go_in;
  wire  invoke19_go_out;
  wire  invoke19_done_in;
  wire  invoke19_done_out;
  wire  invoke20_go_in;
  wire  invoke20_go_out;
  wire  invoke20_done_in;
  wire  invoke20_done_out;
  wire  invoke21_go_in;
  wire  invoke21_go_out;
  wire  invoke21_done_in;
  wire  invoke21_done_out;
  wire  invoke22_go_in;
  wire  invoke22_go_out;
  wire  invoke22_done_in;
  wire  invoke22_done_out;
  wire  invoke23_go_in;
  wire  invoke23_go_out;
  wire  invoke23_done_in;
  wire  invoke23_done_out;
  wire  invoke33_go_in;
  wire  invoke33_go_out;
  wire  invoke33_done_in;
  wire  invoke33_done_out;
  wire  early_reset_cond00_go_in;
  wire  early_reset_cond00_go_out;
  wire  early_reset_cond00_done_in;
  wire  early_reset_cond00_done_out;
  wire  early_reset_cond10_go_in;
  wire  early_reset_cond10_go_out;
  wire  early_reset_cond10_done_in;
  wire  early_reset_cond10_done_out;
  wire  early_reset_cond20_go_in;
  wire  early_reset_cond20_go_out;
  wire  early_reset_cond20_done_in;
  wire  early_reset_cond20_done_out;
  wire  early_reset_static_par_go_in;
  wire  early_reset_static_par_go_out;
  wire  early_reset_static_par_done_in;
  wire  early_reset_static_par_done_out;
  wire  early_reset_static_par0_go_in;
  wire  early_reset_static_par0_go_out;
  wire  early_reset_static_par0_done_in;
  wire  early_reset_static_par0_done_out;
  wire  early_reset_static_seq_go_in;
  wire  early_reset_static_seq_go_out;
  wire  early_reset_static_seq_done_in;
  wire  early_reset_static_seq_done_out;
  wire  early_reset_static_par1_go_in;
  wire  early_reset_static_par1_go_out;
  wire  early_reset_static_par1_done_in;
  wire  early_reset_static_par1_done_out;
  wire  early_reset_static_seq1_go_in;
  wire  early_reset_static_seq1_go_out;
  wire  early_reset_static_seq1_done_in;
  wire  early_reset_static_seq1_done_out;
  wire  wrapper_early_reset_static_par_go_in;
  wire  wrapper_early_reset_static_par_go_out;
  wire  wrapper_early_reset_static_par_done_in;
  wire  wrapper_early_reset_static_par_done_out;
  wire  wrapper_early_reset_cond00_go_in;
  wire  wrapper_early_reset_cond00_go_out;
  wire  wrapper_early_reset_cond00_done_in;
  wire  wrapper_early_reset_cond00_done_out;
  wire  wrapper_early_reset_cond10_go_in;
  wire  wrapper_early_reset_cond10_go_out;
  wire  wrapper_early_reset_cond10_done_in;
  wire  wrapper_early_reset_cond10_done_out;
  wire  wrapper_early_reset_static_par0_go_in;
  wire  wrapper_early_reset_static_par0_go_out;
  wire  wrapper_early_reset_static_par0_done_in;
  wire  wrapper_early_reset_static_par0_done_out;
  wire  wrapper_early_reset_cond20_go_in;
  wire  wrapper_early_reset_cond20_go_out;
  wire  wrapper_early_reset_cond20_done_in;
  wire  wrapper_early_reset_cond20_done_out;
  wire  wrapper_early_reset_static_seq_go_in;
  wire  wrapper_early_reset_static_seq_go_out;
  wire  wrapper_early_reset_static_seq_done_in;
  wire  wrapper_early_reset_static_seq_done_out;
  wire  wrapper_early_reset_static_par1_go_in;
  wire  wrapper_early_reset_static_par1_go_out;
  wire  wrapper_early_reset_static_par1_done_in;
  wire  wrapper_early_reset_static_par1_done_out;
  wire  wrapper_early_reset_static_seq1_go_in;
  wire  wrapper_early_reset_static_seq1_go_out;
  wire  wrapper_early_reset_static_seq1_done_in;
  wire  wrapper_early_reset_static_seq1_done_out;
  wire  par0_go_in;
  wire  par0_go_out;
  wire  par0_done_in;
  wire  par0_done_out;
  wire  tdcc_go_in;
  wire  tdcc_go_out;
  wire  tdcc_done_in;
  wire  tdcc_done_out;
  wire  tdcc0_go_in;
  wire  tdcc0_go_out;
  wire  tdcc0_done_in;
  wire  tdcc0_done_out;
  wire  tdcc1_go_in;
  wire  tdcc1_go_out;
  wire  tdcc1_done_in;
  wire  tdcc1_done_out;
  wire  par1_go_in;
  wire  par1_go_out;
  wire  par1_done_in;
  wire  par1_done_out;
  wire  tdcc2_go_in;
  wire  tdcc2_go_out;
  wire  tdcc2_done_in;
  wire  tdcc2_done_out;
  wire  tdcc3_go_in;
  wire  tdcc3_go_out;
  wire  tdcc3_done_in;
  wire  tdcc3_done_out;
  wire  par2_go_in;
  wire  par2_go_out;
  wire  par2_done_in;
  wire  par2_done_out;
  wire  tdcc4_go_in;
  wire  tdcc4_go_out;
  wire  tdcc4_done_in;
  wire  tdcc4_done_out;
  wire  tdcc5_go_in;
  wire  tdcc5_go_out;
  wire  tdcc5_done_in;
  wire  tdcc5_done_out;
  wire  tdcc6_go_in;
  wire  tdcc6_go_out;
  wire  tdcc6_done_in;
  wire  tdcc6_done_out;
  wire  tdcc7_go_in;
  wire  tdcc7_go_out;
  wire  tdcc7_done_in;
  wire  tdcc7_done_out;
  wire  tdcc8_go_in;
  wire  tdcc8_go_out;
  wire  tdcc8_done_in;
  wire  tdcc8_done_out;
  wire [3:0] _GEN_1 = invoke33_go_out ? add2_out : 4'h0; // @[]
  wire  _GEN_4 = early_reset_cond20_go_out; // @[]
  wire [3:0] _GEN_13 = beg_spl_let17_go_out ? i0_out : 4'h0; // @[]
  wire [31:0] _GEN_15 = fsm_out == 5'h8 & early_reset_static_seq_go_out ? add3_out : 32'h0; // @[]
  wire [3:0] _GEN_17 = beg_spl_let13_go_out | fsm_out == 5'h10 & early_reset_static_seq1_go_out ? i0_out : 4'h0; // @[]
  wire [3:0] _GEN_22 = beg_spl_let16_go_out | beg_spl_let6_go_out ? i0_out : 4'h0; // @[]
  wire [4:0] _GEN_30 = fsm_out != 5'h0 & early_reset_cond20_go_out ? adder1_out : 5'h0; // @[]
  wire [4:0] _GEN_31 = fsm_out != 5'h0 & early_reset_cond00_go_out ? adder_out : _GEN_30; // @[]
  wire [4:0] _GEN_32 = fsm_out != 5'h8 & early_reset_static_seq_go_out ? adder4_out : _GEN_31; // @[]
  wire [4:0] _GEN_33 = fsm_out == 5'h0 & early_reset_cond00_go_out | fsm_out == 5'h0 & early_reset_cond10_go_out |
    fsm_out == 5'h0 & early_reset_cond20_go_out | fsm_out == 5'h0 & early_reset_static_par_go_out | fsm_out == 5'h0 &
    early_reset_static_par0_go_out | fsm_out == 5'h8 & early_reset_static_seq_go_out | fsm_out == 5'h4 &
    early_reset_static_par1_go_out | fsm_out == 5'h11 & early_reset_static_seq1_go_out ? 5'h0 : _GEN_32; // @[]
  wire [4:0] _GEN_34 = fsm_out != 5'h11 & early_reset_static_seq1_go_out ? adder6_out : _GEN_33; // @[]
  wire [4:0] _GEN_35 = fsm_out != 5'h0 & early_reset_static_par_go_out ? adder2_out : _GEN_34; // @[]
  wire [4:0] _GEN_36 = fsm_out != 5'h0 & early_reset_static_par0_go_out ? adder3_out : _GEN_35; // @[]
  wire [4:0] _GEN_37 = fsm_out != 5'h4 & early_reset_static_par1_go_out ? adder5_out : _GEN_36; // @[]
  wire  _GEN_40 = early_reset_cond00_go_out; // @[]
  wire  _GEN_43 = fsm6_out == 2'h2 ? 1'h0 : fsm6_out == 2'h0 & beg_spl_let15_done_out & tdcc5_go_out; // @[]
  wire  _GEN_52 = early_reset_static_seq_go_out; // @[]
  wire  _GEN_55 = fsm3_out == 2'h2 ? 1'h0 : fsm3_out == 2'h0 & beg_spl_let10_done_out & tdcc2_go_out; // @[]
  wire  _GEN_59 = fsm5_out == 2'h2 ? 1'h0 : fsm5_out == 2'h0 & beg_spl_let14_done_out & tdcc4_go_out; // @[]
  wire [31:0] _GEN_68 = invoke8_go_out | invoke14_go_out | invoke23_go_out ? A_int_read_data : 32'h0; // @[]
  wire [3:0] _GEN_70 = invoke33_go_out ? i0_out : 4'h0; // @[]
  wire [3:0] _GEN_71 = fsm_out == 5'h0 & early_reset_static_par1_go_out ? k_0_out : _GEN_70; // @[]
  wire  _GEN_77 = fsm8_out == 2'h2 ? 1'h0 : fsm8_out == 2'h0 & beg_spl_let17_done_out & tdcc7_go_out; // @[]
  wire [31:0] _GEN_80 = fsm_out == 5'h8 & early_reset_static_seq_go_out ? A_int_read0_0_out : 32'h0; // @[]
  wire [31:0] _GEN_81 = fsm_out == 5'h4 & early_reset_static_par1_go_out ? temp2_0_out : _GEN_80; // @[]
  wire [31:0] _GEN_83 = fsm_out == 5'h4 & early_reset_static_par1_go_out | fsm_out == 5'h10 &
    early_reset_static_seq1_go_out ? A_int_read0_0_out : 32'h0; // @[]
  wire  _GEN_91 = fsm1_out == 2'h2 ? 1'h0 : fsm1_out == 2'h0 & beg_spl_let6_done_out & tdcc0_go_out; // @[]
  wire  _GEN_95 = fsm4_out == 2'h2 ? 1'h0 : fsm4_out == 2'h0 & beg_spl_let11_done_out & tdcc3_go_out; // @[]
  wire  _GEN_447 = fsm9_out == 5'h0 & wrapper_early_reset_static_par_done_out & tdcc8_go_out; // @[]
  wire  _GEN_475 = fsm9_out == 5'h4 & wrapper_early_reset_static_par0_done_out & tdcc8_go_out; // @[]
  wire  _GEN_479 = fsm9_out == 5'h14 | fsm9_out == 5'h0 & wrapper_early_reset_static_par_done_out & tdcc8_go_out |
    fsm9_out == 5'h1 & (wrapper_early_reset_cond00_done_out & comb_reg_out) & tdcc8_go_out | fsm9_out == 5'h13 & (
    wrapper_early_reset_cond00_done_out & comb_reg_out) & tdcc8_go_out | fsm9_out == 5'h2 & invoke2_done_out &
    tdcc8_go_out | fsm9_out == 5'h3 & (wrapper_early_reset_cond10_done_out & comb_reg0_out) & tdcc8_go_out | fsm9_out
     == 5'h11 & (wrapper_early_reset_cond10_done_out & comb_reg0_out) & tdcc8_go_out | _GEN_475; // @[]
  wire  _GEN_508 = _GEN_479 | fsm9_out == 5'h5 & (wrapper_early_reset_cond20_done_out & comb_reg1_out) & tdcc8_go_out |
    fsm9_out == 5'hc & (wrapper_early_reset_cond20_done_out & comb_reg1_out) & tdcc8_go_out | fsm9_out == 5'h6 &
    beg_spl_let4_done_out & tdcc8_go_out | fsm9_out == 5'h7 & invoke5_done_out & tdcc8_go_out | fsm9_out == 5'h8 &
    par0_done_out & tdcc8_go_out | fsm9_out == 5'h9 & wrapper_early_reset_static_seq_done_out & tdcc8_go_out | fsm9_out
     == 5'ha & par1_done_out & tdcc8_go_out; // @[]
  wire  _GEN_537 = fsm9_out == 5'h10 & wrapper_early_reset_static_seq1_done_out & tdcc8_go_out; // @[]
  wire  _GEN_543 = fsm9_out == 5'h3 & (wrapper_early_reset_cond10_done_out & ~comb_reg0_out) & tdcc8_go_out; // @[]
  wire  _GEN_548 = _GEN_508 | fsm9_out == 5'hb & wrapper_early_reset_static_par1_done_out & tdcc8_go_out | fsm9_out == 5'h5
     & (wrapper_early_reset_cond20_done_out & ~comb_reg1_out) & tdcc8_go_out | fsm9_out == 5'hc & (
    wrapper_early_reset_cond20_done_out & ~comb_reg1_out) & tdcc8_go_out | fsm9_out == 5'hd & beg_spl_let13_done_out &
    tdcc8_go_out | fsm9_out == 5'he & invoke19_done_out & tdcc8_go_out | fsm9_out == 5'hf & par2_done_out & tdcc8_go_out
     | _GEN_537 | _GEN_543; // @[]
  wire [3:0] _GEN_102 = fsm9_out == 5'he & invoke19_done_out & tdcc8_go_out ? 4'hf : {{3'd0}, _GEN_447}; // @[]
  wire [4:0] _GEN_103 = fsm9_out == 5'h3 & (wrapper_early_reset_cond10_done_out & ~comb_reg0_out) & tdcc8_go_out |
    fsm9_out == 5'h11 & (wrapper_early_reset_cond10_done_out & ~comb_reg0_out) & tdcc8_go_out ? 5'h12 : {{1'd0},
    _GEN_102}; // @[]
  wire [4:0] _GEN_104 = fsm9_out == 5'hf & par2_done_out & tdcc8_go_out ? 5'h10 : _GEN_103; // @[]
  wire [4:0] _GEN_105 = fsm9_out == 5'h14 ? 5'h0 : _GEN_104; // @[]
  wire [4:0] _GEN_106 = fsm9_out == 5'h2 & invoke2_done_out & tdcc8_go_out ? 5'h3 : _GEN_105; // @[]
  wire [4:0] _GEN_107 = fsm9_out == 5'h5 & (wrapper_early_reset_cond20_done_out & ~comb_reg1_out) & tdcc8_go_out |
    fsm9_out == 5'hc & (wrapper_early_reset_cond20_done_out & ~comb_reg1_out) & tdcc8_go_out ? 5'hd : _GEN_106; // @[]
  wire [4:0] _GEN_108 = fsm9_out == 5'hd & beg_spl_let13_done_out & tdcc8_go_out ? 5'he : _GEN_107; // @[]
  wire [4:0] _GEN_109 = fsm9_out == 5'hb & wrapper_early_reset_static_par1_done_out & tdcc8_go_out ? 5'hc : _GEN_108; // @[]
  wire [4:0] _GEN_110 = fsm9_out == 5'h4 & wrapper_early_reset_static_par0_done_out & tdcc8_go_out ? 5'h5 : _GEN_109; // @[]
  wire [4:0] _GEN_111 = fsm9_out == 5'h1 & (wrapper_early_reset_cond00_done_out & comb_reg_out) & tdcc8_go_out |
    fsm9_out == 5'h13 & (wrapper_early_reset_cond00_done_out & comb_reg_out) & tdcc8_go_out ? 5'h2 : _GEN_110; // @[]
  wire [4:0] _GEN_112 = fsm9_out == 5'h7 & invoke5_done_out & tdcc8_go_out ? 5'h8 : _GEN_111; // @[]
  wire [4:0] _GEN_113 = fsm9_out == 5'h9 & wrapper_early_reset_static_seq_done_out & tdcc8_go_out ? 5'ha : _GEN_112; // @[]
  wire [4:0] _GEN_114 = fsm9_out == 5'h6 & beg_spl_let4_done_out & tdcc8_go_out ? 5'h7 : _GEN_113; // @[]
  wire [4:0] _GEN_115 = fsm9_out == 5'ha & par1_done_out & tdcc8_go_out ? 5'hb : _GEN_114; // @[]
  wire [4:0] _GEN_116 = fsm9_out == 5'h12 & invoke33_done_out & tdcc8_go_out ? 5'h13 : _GEN_115; // @[]
  wire [4:0] _GEN_117 = fsm9_out == 5'h3 & (wrapper_early_reset_cond10_done_out & comb_reg0_out) & tdcc8_go_out |
    fsm9_out == 5'h11 & (wrapper_early_reset_cond10_done_out & comb_reg0_out) & tdcc8_go_out ? 5'h4 : _GEN_116; // @[]
  wire [4:0] _GEN_118 = fsm9_out == 5'h1 & (wrapper_early_reset_cond00_done_out & ~comb_reg_out) & tdcc8_go_out |
    fsm9_out == 5'h13 & (wrapper_early_reset_cond00_done_out & ~comb_reg_out) & tdcc8_go_out ? 5'h14 : _GEN_117; // @[]
  wire [4:0] _GEN_119 = fsm9_out == 5'h5 & (wrapper_early_reset_cond20_done_out & comb_reg1_out) & tdcc8_go_out |
    fsm9_out == 5'hc & (wrapper_early_reset_cond20_done_out & comb_reg1_out) & tdcc8_go_out ? 5'h6 : _GEN_118; // @[]
  wire [4:0] _GEN_120 = fsm9_out == 5'h10 & wrapper_early_reset_static_seq1_done_out & tdcc8_go_out ? 5'h11 : _GEN_119; // @[]
  wire [3:0] _GEN_131 = fsm_out == 5'h0 & early_reset_static_par1_go_out ? add2_out : 4'h0; // @[]
  wire  _GEN_133 = early_reset_cond10_go_out; // @[]
  wire  _GEN_136 = early_reset_static_seq1_go_out; // @[]
  wire  _GEN_142 = fsm7_out == 2'h2 ? 1'h0 : fsm7_out == 2'h0 & beg_spl_let16_done_out & tdcc6_go_out; // @[]
  wire  _GEN_149 = early_reset_static_par_go_out; // @[]
  wire  _GEN_152 = fsm0_out == 2'h2 ? 1'h0 : fsm0_out == 2'h0 & beg_spl_let5_done_out & tdcc_go_out; // @[]
  wire  _GEN_156 = fsm2_out == 2'h2 ? 1'h0 : fsm2_out == 2'h0 & beg_spl_let7_done_out & tdcc1_go_out; // @[]
  wire  _GEN_162 = early_reset_static_par0_go_out; // @[]
  wire  _GEN_164 = early_reset_static_par1_go_out; // @[]
  wire [31:0] _GEN_169 = fsm_out < 5'h3 & early_reset_static_seq1_go_out ? beta_int_read0_0_out : 32'h0; // @[]
  wire [31:0] _GEN_170 = fsm_out < 5'h3 & early_reset_static_seq_go_out | (fsm_out >= 5'h4 & fsm_out < 5'h7 | fsm_out
     >= 5'hc & fsm_out < 5'hf) & early_reset_static_seq1_go_out ? alpha_int_read0_0_out : _GEN_169; // @[]
  wire [31:0] _GEN_173 = fsm_out >= 5'h4 & fsm_out < 5'h7 & early_reset_static_seq_go_out | fsm_out < 5'h3 &
    early_reset_static_par1_go_out | fsm_out >= 5'h8 & fsm_out < 5'hb & early_reset_static_seq1_go_out ?
    A_int_read0_0_out : 32'h0; // @[]
  wire [31:0] _GEN_174 = fsm_out >= 5'hc & fsm_out < 5'hf & early_reset_static_seq1_go_out ? temp2_0_out : _GEN_173; // @[]
  wire [31:0] _GEN_175 = fsm_out < 5'h3 & early_reset_static_seq_go_out | fsm_out >= 5'h4 & fsm_out < 5'h7 &
    early_reset_static_seq1_go_out ? B_int_read0_0_out : _GEN_174; // @[]
  wire [31:0] _GEN_178 = early_reset_static_par_go_out | early_reset_static_par0_go_out ? const0_out : 32'h0; // @[]
  wire [3:0] _GEN_188 = early_reset_cond00_go_out ? i0_out : 4'h0; // @[]
  wire [3:0] _GEN_190 = early_reset_cond00_go_out ? const2_out : 4'h0; // @[]
  wire  _GEN_838 = fsm_out == 5'h0 & ~signal_reg_out & wrapper_early_reset_static_seq_go_out; // @[]
  wire  _GEN_843 = fsm_out == 5'h0 & ~signal_reg_out & wrapper_early_reset_static_par1_go_out; // @[]
  wire  _GEN_848 = fsm_out == 5'h0 & ~signal_reg_out & wrapper_early_reset_static_seq1_go_out; // @[]
  wire  _GEN_885 = fsm_out == 5'h0 & ~signal_reg_out & wrapper_early_reset_static_par_go_out | fsm_out == 5'h0 & ~
    signal_reg_out & wrapper_early_reset_cond00_go_out | fsm_out == 5'h0 & ~signal_reg_out &
    wrapper_early_reset_cond10_go_out | fsm_out == 5'h0 & ~signal_reg_out & wrapper_early_reset_static_par0_go_out |
    fsm_out == 5'h0 & ~signal_reg_out & wrapper_early_reset_cond20_go_out | fsm_out == 5'h0 & ~signal_reg_out &
    wrapper_early_reset_static_seq_go_out | _GEN_843; // @[]
  wire [31:0] _GEN_217 = invoke7_go_out | invoke13_go_out | invoke22_go_out ? B_int_read_data : 32'h0; // @[]
  wire [3:0] _GEN_220 = fsm_out == 5'h11 & early_reset_static_seq1_go_out ? add2_out : 4'h0; // @[]
  wire [31:0] _GEN_229 = invoke5_go_out | invoke19_go_out ? C_int_read_data : 32'h0; // @[]
  std_reg #(.WIDTH(32)) A_int_read0_0 (
    .in(A_int_read0_0_in),
    .write_en(A_int_read0_0_write_en),
    .clk(A_int_read0_0_clk),
    .reset(A_int_read0_0_reset),
    .out(A_int_read0_0_out),
    .done(A_int_read0_0_done)
  );
  std_reg #(.WIDTH(32)) B_int_read0_0 (
    .in(B_int_read0_0_in),
    .write_en(B_int_read0_0_write_en),
    .clk(B_int_read0_0_clk),
    .reset(B_int_read0_0_reset),
    .out(B_int_read0_0_out),
    .done(B_int_read0_0_done)
  );
  std_reg #(.WIDTH(32)) C_i_j_0 (
    .in(C_i_j_0_in),
    .write_en(C_i_j_0_write_en),
    .clk(C_i_j_0_clk),
    .reset(C_i_j_0_reset),
    .out(C_i_j_0_out),
    .done(C_i_j_0_done)
  );
  std_add #(.WIDTH(4)) add2 (
    .left(add2_left),
    .right(add2_right),
    .out(add2_out)
  );
  std_add #(.WIDTH(32)) add3 (
    .left(add3_left),
    .right(add3_right),
    .out(add3_out)
  );
  std_add #(.WIDTH(32)) add4 (
    .left(add4_left),
    .right(add4_right),
    .out(add4_out)
  );
  std_reg #(.WIDTH(32)) alpha_int_read0_0 (
    .in(alpha_int_read0_0_in),
    .write_en(alpha_int_read0_0_write_en),
    .clk(alpha_int_read0_0_clk),
    .reset(alpha_int_read0_0_reset),
    .out(alpha_int_read0_0_out),
    .done(alpha_int_read0_0_done)
  );
  std_reg #(.WIDTH(32)) beta_int_read0_0 (
    .in(beta_int_read0_0_in),
    .write_en(beta_int_read0_0_write_en),
    .clk(beta_int_read0_0_clk),
    .reset(beta_int_read0_0_reset),
    .out(beta_int_read0_0_out),
    .done(beta_int_read0_0_done)
  );
  std_const #(.WIDTH(32), .VALUE(0)) const0 (
    .out(const0_out)
  );
  std_const #(.WIDTH(4), .VALUE(0)) const1 (
    .out(const1_out)
  );
  std_const #(.WIDTH(1), .VALUE(0)) const10 (
    .out(const10_out)
  );
  std_const #(.WIDTH(4), .VALUE(1)) const11 (
    .out(const11_out)
  );
  std_const #(.WIDTH(4), .VALUE(7)) const2 (
    .out(const2_out)
  );
  std_const #(.WIDTH(4), .VALUE(11)) const4 (
    .out(const4_out)
  );
  std_const #(.WIDTH(1), .VALUE(0)) const9 (
    .out(const9_out)
  );
  std_reg #(.WIDTH(4)) i0 (
    .in(i0_in),
    .write_en(i0_write_en),
    .clk(i0_clk),
    .reset(i0_reset),
    .out(i0_out),
    .done(i0_done)
  );
  std_reg #(.WIDTH(4)) j0 (
    .in(j0_in),
    .write_en(j0_write_en),
    .clk(j0_clk),
    .reset(j0_reset),
    .out(j0_out),
    .done(j0_done)
  );
  std_reg #(.WIDTH(4)) k_0 (
    .in(k_0_in),
    .write_en(k_0_write_en),
    .clk(k_0_clk),
    .reset(k_0_reset),
    .out(k_0_out),
    .done(k_0_done)
  );
  std_le #(.WIDTH(4)) le0 (
    .left(le0_left),
    .right(le0_right),
    .out(le0_out)
  );
  std_lt #(.WIDTH(4)) lt0 (
    .left(lt0_left),
    .right(lt0_right),
    .out(lt0_out)
  );
  std_mult_pipe #(.WIDTH(32)) mult_pipe0 (
    .clk(mult_pipe0_clk),
    .reset(mult_pipe0_reset),
    .go(mult_pipe0_go),
    .left(mult_pipe0_left),
    .right(mult_pipe0_right),
    .out(mult_pipe0_out),
    .done(mult_pipe0_done)
  );
  std_reg #(.WIDTH(32)) temp2_0 (
    .in(temp2_0_in),
    .write_en(temp2_0_write_en),
    .clk(temp2_0_clk),
    .reset(temp2_0_reset),
    .out(temp2_0_out),
    .done(temp2_0_done)
  );
  std_reg #(.WIDTH(1)) comb_reg (
    .in(comb_reg_in),
    .write_en(comb_reg_write_en),
    .clk(comb_reg_clk),
    .reset(comb_reg_reset),
    .out(comb_reg_out),
    .done(comb_reg_done)
  );
  std_reg #(.WIDTH(1)) comb_reg0 (
    .in(comb_reg0_in),
    .write_en(comb_reg0_write_en),
    .clk(comb_reg0_clk),
    .reset(comb_reg0_reset),
    .out(comb_reg0_out),
    .done(comb_reg0_done)
  );
  std_reg #(.WIDTH(1)) comb_reg1 (
    .in(comb_reg1_in),
    .write_en(comb_reg1_write_en),
    .clk(comb_reg1_clk),
    .reset(comb_reg1_reset),
    .out(comb_reg1_out),
    .done(comb_reg1_done)
  );
  std_reg #(.WIDTH(5)) fsm (
    .in(fsm_in),
    .write_en(fsm_write_en),
    .clk(fsm_clk),
    .reset(fsm_reset),
    .out(fsm_out),
    .done(fsm_done)
  );
  undef #(.WIDTH(1)) ud (
    .out(ud_out)
  );
  std_add #(.WIDTH(5)) adder (
    .left(adder_left),
    .right(adder_right),
    .out(adder_out)
  );
  undef #(.WIDTH(1)) ud0 (
    .out(ud0_out)
  );
  std_add #(.WIDTH(5)) adder0 (
    .left(adder0_left),
    .right(adder0_right),
    .out(adder0_out)
  );
  undef #(.WIDTH(1)) ud1 (
    .out(ud1_out)
  );
  std_add #(.WIDTH(5)) adder1 (
    .left(adder1_left),
    .right(adder1_right),
    .out(adder1_out)
  );
  undef #(.WIDTH(1)) ud2 (
    .out(ud2_out)
  );
  std_add #(.WIDTH(5)) adder2 (
    .left(adder2_left),
    .right(adder2_right),
    .out(adder2_out)
  );
  undef #(.WIDTH(1)) ud3 (
    .out(ud3_out)
  );
  std_add #(.WIDTH(5)) adder3 (
    .left(adder3_left),
    .right(adder3_right),
    .out(adder3_out)
  );
  undef #(.WIDTH(1)) ud4 (
    .out(ud4_out)
  );
  std_add #(.WIDTH(5)) adder4 (
    .left(adder4_left),
    .right(adder4_right),
    .out(adder4_out)
  );
  undef #(.WIDTH(1)) ud5 (
    .out(ud5_out)
  );
  std_add #(.WIDTH(5)) adder5 (
    .left(adder5_left),
    .right(adder5_right),
    .out(adder5_out)
  );
  undef #(.WIDTH(1)) ud6 (
    .out(ud6_out)
  );
  std_add #(.WIDTH(5)) adder6 (
    .left(adder6_left),
    .right(adder6_right),
    .out(adder6_out)
  );
  std_reg #(.WIDTH(1)) signal_reg (
    .in(signal_reg_in),
    .write_en(signal_reg_write_en),
    .clk(signal_reg_clk),
    .reset(signal_reg_reset),
    .out(signal_reg_out),
    .done(signal_reg_done)
  );
  std_reg #(.WIDTH(2)) fsm0 (
    .in(fsm0_in),
    .write_en(fsm0_write_en),
    .clk(fsm0_clk),
    .reset(fsm0_reset),
    .out(fsm0_out),
    .done(fsm0_done)
  );
  std_reg #(.WIDTH(1)) pd (
    .in(pd_in),
    .write_en(pd_write_en),
    .clk(pd_clk),
    .reset(pd_reset),
    .out(pd_out),
    .done(pd_done)
  );
  std_reg #(.WIDTH(2)) fsm1 (
    .in(fsm1_in),
    .write_en(fsm1_write_en),
    .clk(fsm1_clk),
    .reset(fsm1_reset),
    .out(fsm1_out),
    .done(fsm1_done)
  );
  std_reg #(.WIDTH(1)) pd0 (
    .in(pd0_in),
    .write_en(pd0_write_en),
    .clk(pd0_clk),
    .reset(pd0_reset),
    .out(pd0_out),
    .done(pd0_done)
  );
  std_reg #(.WIDTH(2)) fsm2 (
    .in(fsm2_in),
    .write_en(fsm2_write_en),
    .clk(fsm2_clk),
    .reset(fsm2_reset),
    .out(fsm2_out),
    .done(fsm2_done)
  );
  std_reg #(.WIDTH(1)) pd1 (
    .in(pd1_in),
    .write_en(pd1_write_en),
    .clk(pd1_clk),
    .reset(pd1_reset),
    .out(pd1_out),
    .done(pd1_done)
  );
  std_reg #(.WIDTH(2)) fsm3 (
    .in(fsm3_in),
    .write_en(fsm3_write_en),
    .clk(fsm3_clk),
    .reset(fsm3_reset),
    .out(fsm3_out),
    .done(fsm3_done)
  );
  std_reg #(.WIDTH(1)) pd2 (
    .in(pd2_in),
    .write_en(pd2_write_en),
    .clk(pd2_clk),
    .reset(pd2_reset),
    .out(pd2_out),
    .done(pd2_done)
  );
  std_reg #(.WIDTH(2)) fsm4 (
    .in(fsm4_in),
    .write_en(fsm4_write_en),
    .clk(fsm4_clk),
    .reset(fsm4_reset),
    .out(fsm4_out),
    .done(fsm4_done)
  );
  std_reg #(.WIDTH(1)) pd3 (
    .in(pd3_in),
    .write_en(pd3_write_en),
    .clk(pd3_clk),
    .reset(pd3_reset),
    .out(pd3_out),
    .done(pd3_done)
  );
  std_reg #(.WIDTH(2)) fsm5 (
    .in(fsm5_in),
    .write_en(fsm5_write_en),
    .clk(fsm5_clk),
    .reset(fsm5_reset),
    .out(fsm5_out),
    .done(fsm5_done)
  );
  std_reg #(.WIDTH(1)) pd4 (
    .in(pd4_in),
    .write_en(pd4_write_en),
    .clk(pd4_clk),
    .reset(pd4_reset),
    .out(pd4_out),
    .done(pd4_done)
  );
  std_reg #(.WIDTH(2)) fsm6 (
    .in(fsm6_in),
    .write_en(fsm6_write_en),
    .clk(fsm6_clk),
    .reset(fsm6_reset),
    .out(fsm6_out),
    .done(fsm6_done)
  );
  std_reg #(.WIDTH(1)) pd5 (
    .in(pd5_in),
    .write_en(pd5_write_en),
    .clk(pd5_clk),
    .reset(pd5_reset),
    .out(pd5_out),
    .done(pd5_done)
  );
  std_reg #(.WIDTH(2)) fsm7 (
    .in(fsm7_in),
    .write_en(fsm7_write_en),
    .clk(fsm7_clk),
    .reset(fsm7_reset),
    .out(fsm7_out),
    .done(fsm7_done)
  );
  std_reg #(.WIDTH(1)) pd6 (
    .in(pd6_in),
    .write_en(pd6_write_en),
    .clk(pd6_clk),
    .reset(pd6_reset),
    .out(pd6_out),
    .done(pd6_done)
  );
  std_reg #(.WIDTH(2)) fsm8 (
    .in(fsm8_in),
    .write_en(fsm8_write_en),
    .clk(fsm8_clk),
    .reset(fsm8_reset),
    .out(fsm8_out),
    .done(fsm8_done)
  );
  std_reg #(.WIDTH(1)) pd7 (
    .in(pd7_in),
    .write_en(pd7_write_en),
    .clk(pd7_clk),
    .reset(pd7_reset),
    .out(pd7_out),
    .done(pd7_done)
  );
  std_reg #(.WIDTH(5)) fsm9 (
    .in(fsm9_in),
    .write_en(fsm9_write_en),
    .clk(fsm9_clk),
    .reset(fsm9_reset),
    .out(fsm9_out),
    .done(fsm9_done)
  );
  std_wire #(.WIDTH(1)) beg_spl_let10_go (
    .in(beg_spl_let10_go_in),
    .out(beg_spl_let10_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let10_done (
    .in(beg_spl_let10_done_in),
    .out(beg_spl_let10_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let11_go (
    .in(beg_spl_let11_go_in),
    .out(beg_spl_let11_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let11_done (
    .in(beg_spl_let11_done_in),
    .out(beg_spl_let11_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let13_go (
    .in(beg_spl_let13_go_in),
    .out(beg_spl_let13_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let13_done (
    .in(beg_spl_let13_done_in),
    .out(beg_spl_let13_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let14_go (
    .in(beg_spl_let14_go_in),
    .out(beg_spl_let14_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let14_done (
    .in(beg_spl_let14_done_in),
    .out(beg_spl_let14_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let15_go (
    .in(beg_spl_let15_go_in),
    .out(beg_spl_let15_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let15_done (
    .in(beg_spl_let15_done_in),
    .out(beg_spl_let15_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let16_go (
    .in(beg_spl_let16_go_in),
    .out(beg_spl_let16_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let16_done (
    .in(beg_spl_let16_done_in),
    .out(beg_spl_let16_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let17_go (
    .in(beg_spl_let17_go_in),
    .out(beg_spl_let17_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let17_done (
    .in(beg_spl_let17_done_in),
    .out(beg_spl_let17_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let4_go (
    .in(beg_spl_let4_go_in),
    .out(beg_spl_let4_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let4_done (
    .in(beg_spl_let4_done_in),
    .out(beg_spl_let4_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let5_go (
    .in(beg_spl_let5_go_in),
    .out(beg_spl_let5_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let5_done (
    .in(beg_spl_let5_done_in),
    .out(beg_spl_let5_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let6_go (
    .in(beg_spl_let6_go_in),
    .out(beg_spl_let6_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let6_done (
    .in(beg_spl_let6_done_in),
    .out(beg_spl_let6_done_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let7_go (
    .in(beg_spl_let7_go_in),
    .out(beg_spl_let7_go_out)
  );
  std_wire #(.WIDTH(1)) beg_spl_let7_done (
    .in(beg_spl_let7_done_in),
    .out(beg_spl_let7_done_out)
  );
  std_wire #(.WIDTH(1)) invoke2_go (
    .in(invoke2_go_in),
    .out(invoke2_go_out)
  );
  std_wire #(.WIDTH(1)) invoke2_done (
    .in(invoke2_done_in),
    .out(invoke2_done_out)
  );
  std_wire #(.WIDTH(1)) invoke5_go (
    .in(invoke5_go_in),
    .out(invoke5_go_out)
  );
  std_wire #(.WIDTH(1)) invoke5_done (
    .in(invoke5_done_in),
    .out(invoke5_done_out)
  );
  std_wire #(.WIDTH(1)) invoke6_go (
    .in(invoke6_go_in),
    .out(invoke6_go_out)
  );
  std_wire #(.WIDTH(1)) invoke6_done (
    .in(invoke6_done_in),
    .out(invoke6_done_out)
  );
  std_wire #(.WIDTH(1)) invoke7_go (
    .in(invoke7_go_in),
    .out(invoke7_go_out)
  );
  std_wire #(.WIDTH(1)) invoke7_done (
    .in(invoke7_done_in),
    .out(invoke7_done_out)
  );
  std_wire #(.WIDTH(1)) invoke8_go (
    .in(invoke8_go_in),
    .out(invoke8_go_out)
  );
  std_wire #(.WIDTH(1)) invoke8_done (
    .in(invoke8_done_in),
    .out(invoke8_done_out)
  );
  std_wire #(.WIDTH(1)) invoke13_go (
    .in(invoke13_go_in),
    .out(invoke13_go_out)
  );
  std_wire #(.WIDTH(1)) invoke13_done (
    .in(invoke13_done_in),
    .out(invoke13_done_out)
  );
  std_wire #(.WIDTH(1)) invoke14_go (
    .in(invoke14_go_in),
    .out(invoke14_go_out)
  );
  std_wire #(.WIDTH(1)) invoke14_done (
    .in(invoke14_done_in),
    .out(invoke14_done_out)
  );
  std_wire #(.WIDTH(1)) invoke19_go (
    .in(invoke19_go_in),
    .out(invoke19_go_out)
  );
  std_wire #(.WIDTH(1)) invoke19_done (
    .in(invoke19_done_in),
    .out(invoke19_done_out)
  );
  std_wire #(.WIDTH(1)) invoke20_go (
    .in(invoke20_go_in),
    .out(invoke20_go_out)
  );
  std_wire #(.WIDTH(1)) invoke20_done (
    .in(invoke20_done_in),
    .out(invoke20_done_out)
  );
  std_wire #(.WIDTH(1)) invoke21_go (
    .in(invoke21_go_in),
    .out(invoke21_go_out)
  );
  std_wire #(.WIDTH(1)) invoke21_done (
    .in(invoke21_done_in),
    .out(invoke21_done_out)
  );
  std_wire #(.WIDTH(1)) invoke22_go (
    .in(invoke22_go_in),
    .out(invoke22_go_out)
  );
  std_wire #(.WIDTH(1)) invoke22_done (
    .in(invoke22_done_in),
    .out(invoke22_done_out)
  );
  std_wire #(.WIDTH(1)) invoke23_go (
    .in(invoke23_go_in),
    .out(invoke23_go_out)
  );
  std_wire #(.WIDTH(1)) invoke23_done (
    .in(invoke23_done_in),
    .out(invoke23_done_out)
  );
  std_wire #(.WIDTH(1)) invoke33_go (
    .in(invoke33_go_in),
    .out(invoke33_go_out)
  );
  std_wire #(.WIDTH(1)) invoke33_done (
    .in(invoke33_done_in),
    .out(invoke33_done_out)
  );
  std_wire #(.WIDTH(1)) early_reset_cond00_go (
    .in(early_reset_cond00_go_in),
    .out(early_reset_cond00_go_out)
  );
  std_wire #(.WIDTH(1)) early_reset_cond00_done (
    .in(early_reset_cond00_done_in),
    .out(early_reset_cond00_done_out)
  );
  std_wire #(.WIDTH(1)) early_reset_cond10_go (
    .in(early_reset_cond10_go_in),
    .out(early_reset_cond10_go_out)
  );
  std_wire #(.WIDTH(1)) early_reset_cond10_done (
    .in(early_reset_cond10_done_in),
    .out(early_reset_cond10_done_out)
  );
  std_wire #(.WIDTH(1)) early_reset_cond20_go (
    .in(early_reset_cond20_go_in),
    .out(early_reset_cond20_go_out)
  );
  std_wire #(.WIDTH(1)) early_reset_cond20_done (
    .in(early_reset_cond20_done_in),
    .out(early_reset_cond20_done_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_par_go (
    .in(early_reset_static_par_go_in),
    .out(early_reset_static_par_go_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_par_done (
    .in(early_reset_static_par_done_in),
    .out(early_reset_static_par_done_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_par0_go (
    .in(early_reset_static_par0_go_in),
    .out(early_reset_static_par0_go_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_par0_done (
    .in(early_reset_static_par0_done_in),
    .out(early_reset_static_par0_done_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_seq_go (
    .in(early_reset_static_seq_go_in),
    .out(early_reset_static_seq_go_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_seq_done (
    .in(early_reset_static_seq_done_in),
    .out(early_reset_static_seq_done_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_par1_go (
    .in(early_reset_static_par1_go_in),
    .out(early_reset_static_par1_go_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_par1_done (
    .in(early_reset_static_par1_done_in),
    .out(early_reset_static_par1_done_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_seq1_go (
    .in(early_reset_static_seq1_go_in),
    .out(early_reset_static_seq1_go_out)
  );
  std_wire #(.WIDTH(1)) early_reset_static_seq1_done (
    .in(early_reset_static_seq1_done_in),
    .out(early_reset_static_seq1_done_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_par_go (
    .in(wrapper_early_reset_static_par_go_in),
    .out(wrapper_early_reset_static_par_go_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_par_done (
    .in(wrapper_early_reset_static_par_done_in),
    .out(wrapper_early_reset_static_par_done_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_cond00_go (
    .in(wrapper_early_reset_cond00_go_in),
    .out(wrapper_early_reset_cond00_go_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_cond00_done (
    .in(wrapper_early_reset_cond00_done_in),
    .out(wrapper_early_reset_cond00_done_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_cond10_go (
    .in(wrapper_early_reset_cond10_go_in),
    .out(wrapper_early_reset_cond10_go_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_cond10_done (
    .in(wrapper_early_reset_cond10_done_in),
    .out(wrapper_early_reset_cond10_done_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_par0_go (
    .in(wrapper_early_reset_static_par0_go_in),
    .out(wrapper_early_reset_static_par0_go_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_par0_done (
    .in(wrapper_early_reset_static_par0_done_in),
    .out(wrapper_early_reset_static_par0_done_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_cond20_go (
    .in(wrapper_early_reset_cond20_go_in),
    .out(wrapper_early_reset_cond20_go_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_cond20_done (
    .in(wrapper_early_reset_cond20_done_in),
    .out(wrapper_early_reset_cond20_done_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_seq_go (
    .in(wrapper_early_reset_static_seq_go_in),
    .out(wrapper_early_reset_static_seq_go_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_seq_done (
    .in(wrapper_early_reset_static_seq_done_in),
    .out(wrapper_early_reset_static_seq_done_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_par1_go (
    .in(wrapper_early_reset_static_par1_go_in),
    .out(wrapper_early_reset_static_par1_go_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_par1_done (
    .in(wrapper_early_reset_static_par1_done_in),
    .out(wrapper_early_reset_static_par1_done_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_seq1_go (
    .in(wrapper_early_reset_static_seq1_go_in),
    .out(wrapper_early_reset_static_seq1_go_out)
  );
  std_wire #(.WIDTH(1)) wrapper_early_reset_static_seq1_done (
    .in(wrapper_early_reset_static_seq1_done_in),
    .out(wrapper_early_reset_static_seq1_done_out)
  );
  std_wire #(.WIDTH(1)) par0_go (
    .in(par0_go_in),
    .out(par0_go_out)
  );
  std_wire #(.WIDTH(1)) par0_done (
    .in(par0_done_in),
    .out(par0_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc_go (
    .in(tdcc_go_in),
    .out(tdcc_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc_done (
    .in(tdcc_done_in),
    .out(tdcc_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc0_go (
    .in(tdcc0_go_in),
    .out(tdcc0_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc0_done (
    .in(tdcc0_done_in),
    .out(tdcc0_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc1_go (
    .in(tdcc1_go_in),
    .out(tdcc1_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc1_done (
    .in(tdcc1_done_in),
    .out(tdcc1_done_out)
  );
  std_wire #(.WIDTH(1)) par1_go (
    .in(par1_go_in),
    .out(par1_go_out)
  );
  std_wire #(.WIDTH(1)) par1_done (
    .in(par1_done_in),
    .out(par1_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc2_go (
    .in(tdcc2_go_in),
    .out(tdcc2_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc2_done (
    .in(tdcc2_done_in),
    .out(tdcc2_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc3_go (
    .in(tdcc3_go_in),
    .out(tdcc3_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc3_done (
    .in(tdcc3_done_in),
    .out(tdcc3_done_out)
  );
  std_wire #(.WIDTH(1)) par2_go (
    .in(par2_go_in),
    .out(par2_go_out)
  );
  std_wire #(.WIDTH(1)) par2_done (
    .in(par2_done_in),
    .out(par2_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc4_go (
    .in(tdcc4_go_in),
    .out(tdcc4_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc4_done (
    .in(tdcc4_done_in),
    .out(tdcc4_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc5_go (
    .in(tdcc5_go_in),
    .out(tdcc5_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc5_done (
    .in(tdcc5_done_in),
    .out(tdcc5_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc6_go (
    .in(tdcc6_go_in),
    .out(tdcc6_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc6_done (
    .in(tdcc6_done_in),
    .out(tdcc6_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc7_go (
    .in(tdcc7_go_in),
    .out(tdcc7_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc7_done (
    .in(tdcc7_done_in),
    .out(tdcc7_done_out)
  );
  std_wire #(.WIDTH(1)) tdcc8_go (
    .in(tdcc8_go_in),
    .out(tdcc8_go_out)
  );
  std_wire #(.WIDTH(1)) tdcc8_done (
    .in(tdcc8_done_in),
    .out(tdcc8_done_out)
  );
  assign done = tdcc8_done_out; // @[]
  assign A_int_addr0 = beg_spl_let11_go_out | beg_spl_let17_go_out | beg_spl_let7_go_out ? i0_out : 4'h0; // @[]
  assign A_int_addr1 = beg_spl_let11_go_out | beg_spl_let7_go_out ? k_0_out : _GEN_13; // @[]
  assign A_int_write_en = 1'h0;
  assign A_int_write_data = 32'h0;
  assign A_int_read_en = beg_spl_let11_go_out | beg_spl_let17_go_out | beg_spl_let7_go_out; // @[]
  assign B_int_addr0 = beg_spl_let10_go_out ? k_0_out : _GEN_22; // @[]
  assign B_int_addr1 = beg_spl_let10_go_out | beg_spl_let16_go_out | beg_spl_let6_go_out ? j0_out : 4'h0; // @[]
  assign B_int_write_en = 1'h0;
  assign B_int_write_data = 32'h0;
  assign B_int_read_en = beg_spl_let10_go_out | beg_spl_let16_go_out | beg_spl_let6_go_out; // @[]
  assign C_int_addr0 = beg_spl_let4_go_out | fsm_out == 5'h8 & early_reset_static_seq_go_out ? k_0_out : _GEN_17; // @[]
  assign C_int_addr1 = beg_spl_let13_go_out | beg_spl_let4_go_out | fsm_out == 5'h8 & early_reset_static_seq_go_out |
    fsm_out == 5'h10 & early_reset_static_seq1_go_out ? j0_out : 4'h0; // @[]
  assign C_int_write_en = fsm_out == 5'h8 & early_reset_static_seq_go_out | fsm_out == 5'h10 &
    early_reset_static_seq1_go_out; // @[]
  assign C_int_write_data = fsm_out == 5'h10 & early_reset_static_seq1_go_out ? add4_out : _GEN_15; // @[]
  assign C_int_read_en = beg_spl_let13_go_out | beg_spl_let4_go_out; // @[]
  assign alpha_int_addr0 = (beg_spl_let15_go_out | beg_spl_let5_go_out) & const10_out; // @[]
  assign alpha_int_write_en = 1'h0;
  assign alpha_int_write_data = 32'h0;
  assign alpha_int_read_en = beg_spl_let15_go_out | beg_spl_let5_go_out; // @[]
  assign beta_int_addr0 = beg_spl_let14_go_out & const9_out; // @[]
  assign beta_int_write_en = 1'h0;
  assign beta_int_write_data = 32'h0;
  assign beta_int_read_en = beg_spl_let14_go_out; // @[]
  assign A_int_read0_0_in = fsm_out == 5'h7 & early_reset_static_seq_go_out | fsm_out == 5'h3 &
    early_reset_static_par1_go_out | fsm_out == 5'hb & early_reset_static_seq1_go_out ? mult_pipe0_out : _GEN_68; // @[]
  assign A_int_read0_0_write_en = invoke8_go_out | invoke14_go_out | invoke23_go_out | fsm_out == 5'h7 &
    early_reset_static_seq_go_out | fsm_out == 5'h3 & early_reset_static_par1_go_out | fsm_out == 5'hb &
    early_reset_static_seq1_go_out; // @[]
  assign A_int_read0_0_clk = clk;
  assign A_int_read0_0_reset = reset;
  assign B_int_read0_0_in = fsm_out == 5'h3 & early_reset_static_seq_go_out | (fsm_out == 5'h7 | fsm_out == 5'hf) &
    early_reset_static_seq1_go_out ? mult_pipe0_out : _GEN_217; // @[]
  assign B_int_read0_0_write_en = invoke7_go_out | invoke13_go_out | invoke22_go_out | fsm_out == 5'h3 &
    early_reset_static_seq_go_out | (fsm_out == 5'h7 | fsm_out == 5'hf) & early_reset_static_seq1_go_out; // @[]
  assign B_int_read0_0_clk = clk;
  assign B_int_read0_0_reset = reset;
  assign C_i_j_0_in = fsm_out == 5'h3 & early_reset_static_seq1_go_out ? mult_pipe0_out : _GEN_229; // @[]
  assign C_i_j_0_write_en = invoke5_go_out | invoke19_go_out | fsm_out == 5'h3 & early_reset_static_seq1_go_out; // @[]
  assign C_i_j_0_clk = clk;
  assign C_i_j_0_reset = reset;
  assign add2_left = fsm_out == 5'h11 & early_reset_static_seq1_go_out ? j0_out : _GEN_71; // @[]
  assign add2_right = invoke33_go_out | fsm_out == 5'h0 & early_reset_static_par1_go_out | fsm_out == 5'h11 &
    early_reset_static_seq1_go_out ? const11_out : 4'h0; // @[]
  assign add3_left = fsm_out == 5'h10 & early_reset_static_seq1_go_out ? C_i_j_0_out : _GEN_81; // @[]
  assign add3_right = fsm_out == 5'h8 & early_reset_static_seq_go_out ? C_i_j_0_out : _GEN_83; // @[]
  assign add4_left = fsm_out == 5'h10 & early_reset_static_seq1_go_out ? add3_out : 32'h0; // @[]
  assign add4_right = fsm_out == 5'h10 & early_reset_static_seq1_go_out ? B_int_read0_0_out : 32'h0; // @[]
  assign alpha_int_read0_0_in = invoke6_go_out | invoke21_go_out ? alpha_int_read_data : 32'h0; // @[]
  assign alpha_int_read0_0_write_en = invoke6_go_out | invoke21_go_out; // @[]
  assign alpha_int_read0_0_clk = clk;
  assign alpha_int_read0_0_reset = reset;
  assign beta_int_read0_0_in = invoke20_go_out ? beta_int_read_data : 32'h0; // @[]
  assign beta_int_read0_0_write_en = invoke20_go_out; // @[]
  assign beta_int_read0_0_clk = clk;
  assign beta_int_read0_0_reset = reset;
  assign i0_in = early_reset_static_par_go_out ? const1_out : _GEN_1; // @[]
  assign i0_write_en = invoke33_go_out | early_reset_static_par_go_out; // @[]
  assign i0_clk = clk;
  assign i0_reset = reset;
  assign j0_in = invoke2_go_out ? const1_out : _GEN_220; // @[]
  assign j0_write_en = invoke2_go_out | fsm_out == 5'h11 & early_reset_static_seq1_go_out; // @[]
  assign j0_clk = clk;
  assign j0_reset = reset;
  assign k_0_in = early_reset_static_par0_go_out ? const1_out : _GEN_131; // @[]
  assign k_0_write_en = early_reset_static_par0_go_out | fsm_out == 5'h0 & early_reset_static_par1_go_out; // @[]
  assign k_0_clk = clk;
  assign k_0_reset = reset;
  assign le0_left = early_reset_cond10_go_out ? j0_out : _GEN_188; // @[]
  assign le0_right = early_reset_cond10_go_out ? const4_out : _GEN_190; // @[]
  assign lt0_left = early_reset_cond20_go_out ? k_0_out : 4'h0; // @[]
  assign lt0_right = early_reset_cond20_go_out ? i0_out : 4'h0; // @[]
  assign mult_pipe0_clk = clk;
  assign mult_pipe0_reset = reset;
  assign mult_pipe0_go = (fsm_out < 5'h3 | fsm_out >= 5'h4 & fsm_out < 5'h7) & early_reset_static_seq_go_out | fsm_out
     < 5'h3 & early_reset_static_par1_go_out | (fsm_out < 5'h3 | fsm_out >= 5'h4 & fsm_out < 5'h7 | fsm_out >= 5'h8 &
    fsm_out < 5'hb | fsm_out >= 5'hc & fsm_out < 5'hf) & early_reset_static_seq1_go_out; // @[]
  assign mult_pipe0_left = fsm_out >= 5'h4 & fsm_out < 5'h7 & early_reset_static_seq_go_out | fsm_out < 5'h3 &
    early_reset_static_par1_go_out | fsm_out >= 5'h8 & fsm_out < 5'hb & early_reset_static_seq1_go_out ?
    B_int_read0_0_out : _GEN_170; // @[]
  assign mult_pipe0_right = fsm_out < 5'h3 & early_reset_static_seq1_go_out ? C_i_j_0_out : _GEN_175; // @[]
  assign temp2_0_in = fsm_out == 5'h4 & early_reset_static_par1_go_out ? add3_out : _GEN_178; // @[]
  assign temp2_0_write_en = early_reset_static_par_go_out | early_reset_static_par0_go_out | fsm_out == 5'h4 &
    early_reset_static_par1_go_out; // @[]
  assign temp2_0_clk = clk;
  assign temp2_0_reset = reset;
  assign comb_reg_in = early_reset_cond00_go_out & le0_out; // @[]
  assign comb_reg_write_en = early_reset_cond00_go_out; // @[]
  assign comb_reg_clk = clk;
  assign comb_reg_reset = reset;
  assign comb_reg0_in = early_reset_cond10_go_out & le0_out; // @[]
  assign comb_reg0_write_en = early_reset_cond10_go_out; // @[]
  assign comb_reg0_clk = clk;
  assign comb_reg0_reset = reset;
  assign comb_reg1_in = early_reset_cond20_go_out & lt0_out; // @[]
  assign comb_reg1_write_en = early_reset_cond20_go_out; // @[]
  assign comb_reg1_clk = clk;
  assign comb_reg1_reset = reset;
  assign fsm_in = fsm_out != 5'h0 & early_reset_cond10_go_out ? adder0_out : _GEN_37; // @[]
  assign fsm_write_en = early_reset_cond00_go_out | early_reset_cond10_go_out | early_reset_cond20_go_out |
    early_reset_static_par_go_out | early_reset_static_par0_go_out | early_reset_static_seq_go_out |
    early_reset_static_par1_go_out | early_reset_static_seq1_go_out; // @[]
  assign fsm_clk = clk;
  assign fsm_reset = reset;
  assign adder_left = early_reset_cond00_go_out ? fsm_out : 5'h0; // @[]
  assign adder_right = {{4'd0}, _GEN_40};
  assign adder0_left = early_reset_cond10_go_out ? fsm_out : 5'h0; // @[]
  assign adder0_right = {{4'd0}, _GEN_133};
  assign adder1_left = early_reset_cond20_go_out ? fsm_out : 5'h0; // @[]
  assign adder1_right = {{4'd0}, _GEN_4};
  assign adder2_left = early_reset_static_par_go_out ? fsm_out : 5'h0; // @[]
  assign adder2_right = {{4'd0}, _GEN_149};
  assign adder3_left = early_reset_static_par0_go_out ? fsm_out : 5'h0; // @[]
  assign adder3_right = {{4'd0}, _GEN_162};
  assign adder4_left = early_reset_static_seq_go_out ? fsm_out : 5'h0; // @[]
  assign adder4_right = {{4'd0}, _GEN_52};
  assign adder5_left = early_reset_static_par1_go_out ? fsm_out : 5'h0; // @[]
  assign adder5_right = {{4'd0}, _GEN_164};
  assign adder6_left = early_reset_static_seq1_go_out ? fsm_out : 5'h0; // @[]
  assign adder6_right = {{4'd0}, _GEN_136};
  assign signal_reg_in = fsm_out == 5'h0 & signal_reg_out ? 1'h0 : _GEN_885 | fsm_out == 5'h0 & ~signal_reg_out &
    wrapper_early_reset_static_seq1_go_out; // @[]
  assign signal_reg_write_en = fsm_out == 5'h0 & signal_reg_out | fsm_out == 5'h0 & ~signal_reg_out &
    wrapper_early_reset_static_par_go_out | fsm_out == 5'h0 & ~signal_reg_out & wrapper_early_reset_cond00_go_out |
    fsm_out == 5'h0 & ~signal_reg_out & wrapper_early_reset_cond10_go_out | fsm_out == 5'h0 & ~signal_reg_out &
    wrapper_early_reset_static_par0_go_out | fsm_out == 5'h0 & ~signal_reg_out & wrapper_early_reset_cond20_go_out |
    _GEN_838 | _GEN_843 | _GEN_848; // @[]
  assign signal_reg_clk = clk;
  assign signal_reg_reset = reset;
  assign fsm0_in = fsm0_out == 2'h1 & invoke6_done_out & tdcc_go_out ? 2'h2 : {{1'd0}, _GEN_152}; // @[]
  assign fsm0_write_en = fsm0_out == 2'h2 | fsm0_out == 2'h0 & beg_spl_let5_done_out & tdcc_go_out | fsm0_out == 2'h1 &
    invoke6_done_out & tdcc_go_out; // @[]
  assign fsm0_clk = clk;
  assign fsm0_reset = reset;
  assign pd_in = pd_out & pd0_out & pd1_out ? 1'h0 : tdcc_done_out & par0_go_out; // @[]
  assign pd_write_en = pd_out & pd0_out & pd1_out | tdcc_done_out & par0_go_out; // @[]
  assign pd_clk = clk;
  assign pd_reset = reset;
  assign fsm1_in = fsm1_out == 2'h1 & invoke7_done_out & tdcc0_go_out ? 2'h2 : {{1'd0}, _GEN_91}; // @[]
  assign fsm1_write_en = fsm1_out == 2'h2 | fsm1_out == 2'h0 & beg_spl_let6_done_out & tdcc0_go_out | fsm1_out == 2'h1
     & invoke7_done_out & tdcc0_go_out; // @[]
  assign fsm1_clk = clk;
  assign fsm1_reset = reset;
  assign pd0_in = pd_out & pd0_out & pd1_out ? 1'h0 : tdcc0_done_out & par0_go_out; // @[]
  assign pd0_write_en = pd_out & pd0_out & pd1_out | tdcc0_done_out & par0_go_out; // @[]
  assign pd0_clk = clk;
  assign pd0_reset = reset;
  assign fsm2_in = fsm2_out == 2'h1 & invoke8_done_out & tdcc1_go_out ? 2'h2 : {{1'd0}, _GEN_156}; // @[]
  assign fsm2_write_en = fsm2_out == 2'h2 | fsm2_out == 2'h0 & beg_spl_let7_done_out & tdcc1_go_out | fsm2_out == 2'h1
     & invoke8_done_out & tdcc1_go_out; // @[]
  assign fsm2_clk = clk;
  assign fsm2_reset = reset;
  assign pd1_in = pd_out & pd0_out & pd1_out ? 1'h0 : tdcc1_done_out & par0_go_out; // @[]
  assign pd1_write_en = pd_out & pd0_out & pd1_out | tdcc1_done_out & par0_go_out; // @[]
  assign pd1_clk = clk;
  assign pd1_reset = reset;
  assign fsm3_in = fsm3_out == 2'h1 & invoke13_done_out & tdcc2_go_out ? 2'h2 : {{1'd0}, _GEN_55}; // @[]
  assign fsm3_write_en = fsm3_out == 2'h2 | fsm3_out == 2'h0 & beg_spl_let10_done_out & tdcc2_go_out | fsm3_out == 2'h1
     & invoke13_done_out & tdcc2_go_out; // @[]
  assign fsm3_clk = clk;
  assign fsm3_reset = reset;
  assign pd2_in = pd2_out & pd3_out ? 1'h0 : tdcc2_done_out & par1_go_out; // @[]
  assign pd2_write_en = pd2_out & pd3_out | tdcc2_done_out & par1_go_out; // @[]
  assign pd2_clk = clk;
  assign pd2_reset = reset;
  assign fsm4_in = fsm4_out == 2'h1 & invoke14_done_out & tdcc3_go_out ? 2'h2 : {{1'd0}, _GEN_95}; // @[]
  assign fsm4_write_en = fsm4_out == 2'h2 | fsm4_out == 2'h0 & beg_spl_let11_done_out & tdcc3_go_out | fsm4_out == 2'h1
     & invoke14_done_out & tdcc3_go_out; // @[]
  assign fsm4_clk = clk;
  assign fsm4_reset = reset;
  assign pd3_in = pd2_out & pd3_out ? 1'h0 : tdcc3_done_out & par1_go_out; // @[]
  assign pd3_write_en = pd2_out & pd3_out | tdcc3_done_out & par1_go_out; // @[]
  assign pd3_clk = clk;
  assign pd3_reset = reset;
  assign fsm5_in = fsm5_out == 2'h1 & invoke20_done_out & tdcc4_go_out ? 2'h2 : {{1'd0}, _GEN_59}; // @[]
  assign fsm5_write_en = fsm5_out == 2'h2 | fsm5_out == 2'h0 & beg_spl_let14_done_out & tdcc4_go_out | fsm5_out == 2'h1
     & invoke20_done_out & tdcc4_go_out; // @[]
  assign fsm5_clk = clk;
  assign fsm5_reset = reset;
  assign pd4_in = pd4_out & pd5_out & pd6_out & pd7_out ? 1'h0 : tdcc4_done_out & par2_go_out; // @[]
  assign pd4_write_en = pd4_out & pd5_out & pd6_out & pd7_out | tdcc4_done_out & par2_go_out; // @[]
  assign pd4_clk = clk;
  assign pd4_reset = reset;
  assign fsm6_in = fsm6_out == 2'h1 & invoke21_done_out & tdcc5_go_out ? 2'h2 : {{1'd0}, _GEN_43}; // @[]
  assign fsm6_write_en = fsm6_out == 2'h2 | fsm6_out == 2'h0 & beg_spl_let15_done_out & tdcc5_go_out | fsm6_out == 2'h1
     & invoke21_done_out & tdcc5_go_out; // @[]
  assign fsm6_clk = clk;
  assign fsm6_reset = reset;
  assign pd5_in = pd4_out & pd5_out & pd6_out & pd7_out ? 1'h0 : tdcc5_done_out & par2_go_out; // @[]
  assign pd5_write_en = pd4_out & pd5_out & pd6_out & pd7_out | tdcc5_done_out & par2_go_out; // @[]
  assign pd5_clk = clk;
  assign pd5_reset = reset;
  assign fsm7_in = fsm7_out == 2'h1 & invoke22_done_out & tdcc6_go_out ? 2'h2 : {{1'd0}, _GEN_142}; // @[]
  assign fsm7_write_en = fsm7_out == 2'h2 | fsm7_out == 2'h0 & beg_spl_let16_done_out & tdcc6_go_out | fsm7_out == 2'h1
     & invoke22_done_out & tdcc6_go_out; // @[]
  assign fsm7_clk = clk;
  assign fsm7_reset = reset;
  assign pd6_in = pd4_out & pd5_out & pd6_out & pd7_out ? 1'h0 : tdcc6_done_out & par2_go_out; // @[]
  assign pd6_write_en = pd4_out & pd5_out & pd6_out & pd7_out | tdcc6_done_out & par2_go_out; // @[]
  assign pd6_clk = clk;
  assign pd6_reset = reset;
  assign fsm8_in = fsm8_out == 2'h1 & invoke23_done_out & tdcc7_go_out ? 2'h2 : {{1'd0}, _GEN_77}; // @[]
  assign fsm8_write_en = fsm8_out == 2'h2 | fsm8_out == 2'h0 & beg_spl_let17_done_out & tdcc7_go_out | fsm8_out == 2'h1
     & invoke23_done_out & tdcc7_go_out; // @[]
  assign fsm8_clk = clk;
  assign fsm8_reset = reset;
  assign pd7_in = pd4_out & pd5_out & pd6_out & pd7_out ? 1'h0 : tdcc7_done_out & par2_go_out; // @[]
  assign pd7_write_en = pd4_out & pd5_out & pd6_out & pd7_out | tdcc7_done_out & par2_go_out; // @[]
  assign pd7_clk = clk;
  assign pd7_reset = reset;
  assign fsm9_in = fsm9_out == 5'h8 & par0_done_out & tdcc8_go_out ? 5'h9 : _GEN_120; // @[]
  assign fsm9_write_en = _GEN_548 | fsm9_out == 5'h11 & (wrapper_early_reset_cond10_done_out & ~comb_reg0_out) &
    tdcc8_go_out | fsm9_out == 5'h12 & invoke33_done_out & tdcc8_go_out | fsm9_out == 5'h1 & (
    wrapper_early_reset_cond00_done_out & ~comb_reg_out) & tdcc8_go_out | fsm9_out == 5'h13 & (
    wrapper_early_reset_cond00_done_out & ~comb_reg_out) & tdcc8_go_out; // @[]
  assign fsm9_clk = clk;
  assign fsm9_reset = reset;
  assign beg_spl_let10_go_in = ~beg_spl_let10_done_out & fsm3_out == 2'h0 & tdcc2_go_out; // @[]
  assign beg_spl_let10_done_in = B_int_read_done;
  assign beg_spl_let11_go_in = ~beg_spl_let11_done_out & fsm4_out == 2'h0 & tdcc3_go_out; // @[]
  assign beg_spl_let11_done_in = A_int_read_done;
  assign beg_spl_let13_go_in = ~beg_spl_let13_done_out & fsm9_out == 5'hd & tdcc8_go_out; // @[]
  assign beg_spl_let13_done_in = C_int_read_done;
  assign beg_spl_let14_go_in = ~beg_spl_let14_done_out & fsm5_out == 2'h0 & tdcc4_go_out; // @[]
  assign beg_spl_let14_done_in = beta_int_read_done;
  assign beg_spl_let15_go_in = ~beg_spl_let15_done_out & fsm6_out == 2'h0 & tdcc5_go_out; // @[]
  assign beg_spl_let15_done_in = alpha_int_read_done;
  assign beg_spl_let16_go_in = ~beg_spl_let16_done_out & fsm7_out == 2'h0 & tdcc6_go_out; // @[]
  assign beg_spl_let16_done_in = B_int_read_done;
  assign beg_spl_let17_go_in = ~beg_spl_let17_done_out & fsm8_out == 2'h0 & tdcc7_go_out; // @[]
  assign beg_spl_let17_done_in = A_int_read_done;
  assign beg_spl_let4_go_in = ~beg_spl_let4_done_out & fsm9_out == 5'h6 & tdcc8_go_out; // @[]
  assign beg_spl_let4_done_in = C_int_read_done;
  assign beg_spl_let5_go_in = ~beg_spl_let5_done_out & fsm0_out == 2'h0 & tdcc_go_out; // @[]
  assign beg_spl_let5_done_in = alpha_int_read_done;
  assign beg_spl_let6_go_in = ~beg_spl_let6_done_out & fsm1_out == 2'h0 & tdcc0_go_out; // @[]
  assign beg_spl_let6_done_in = B_int_read_done;
  assign beg_spl_let7_go_in = ~beg_spl_let7_done_out & fsm2_out == 2'h0 & tdcc1_go_out; // @[]
  assign beg_spl_let7_done_in = A_int_read_done;
  assign invoke2_go_in = ~invoke2_done_out & fsm9_out == 5'h2 & tdcc8_go_out; // @[]
  assign invoke2_done_in = j0_done;
  assign invoke5_go_in = ~invoke5_done_out & fsm9_out == 5'h7 & tdcc8_go_out; // @[]
  assign invoke5_done_in = C_i_j_0_done;
  assign invoke6_go_in = ~invoke6_done_out & fsm0_out == 2'h1 & tdcc_go_out; // @[]
  assign invoke6_done_in = alpha_int_read0_0_done;
  assign invoke7_go_in = ~invoke7_done_out & fsm1_out == 2'h1 & tdcc0_go_out; // @[]
  assign invoke7_done_in = B_int_read0_0_done;
  assign invoke8_go_in = ~invoke8_done_out & fsm2_out == 2'h1 & tdcc1_go_out; // @[]
  assign invoke8_done_in = A_int_read0_0_done;
  assign invoke13_go_in = ~invoke13_done_out & fsm3_out == 2'h1 & tdcc2_go_out; // @[]
  assign invoke13_done_in = B_int_read0_0_done;
  assign invoke14_go_in = ~invoke14_done_out & fsm4_out == 2'h1 & tdcc3_go_out; // @[]
  assign invoke14_done_in = A_int_read0_0_done;
  assign invoke19_go_in = ~invoke19_done_out & fsm9_out == 5'he & tdcc8_go_out; // @[]
  assign invoke19_done_in = C_i_j_0_done;
  assign invoke20_go_in = ~invoke20_done_out & fsm5_out == 2'h1 & tdcc4_go_out; // @[]
  assign invoke20_done_in = beta_int_read0_0_done;
  assign invoke21_go_in = ~invoke21_done_out & fsm6_out == 2'h1 & tdcc5_go_out; // @[]
  assign invoke21_done_in = alpha_int_read0_0_done;
  assign invoke22_go_in = ~invoke22_done_out & fsm7_out == 2'h1 & tdcc6_go_out; // @[]
  assign invoke22_done_in = B_int_read0_0_done;
  assign invoke23_go_in = ~invoke23_done_out & fsm8_out == 2'h1 & tdcc7_go_out; // @[]
  assign invoke23_done_in = A_int_read0_0_done;
  assign invoke33_go_in = ~invoke33_done_out & fsm9_out == 5'h12 & tdcc8_go_out; // @[]
  assign invoke33_done_in = i0_done;
  assign early_reset_cond00_go_in = wrapper_early_reset_cond00_go_out; // @[]
  assign early_reset_cond00_done_in = ud_out;
  assign early_reset_cond10_go_in = wrapper_early_reset_cond10_go_out; // @[]
  assign early_reset_cond10_done_in = ud0_out;
  assign early_reset_cond20_go_in = wrapper_early_reset_cond20_go_out; // @[]
  assign early_reset_cond20_done_in = ud1_out;
  assign early_reset_static_par_go_in = wrapper_early_reset_static_par_go_out; // @[]
  assign early_reset_static_par_done_in = ud2_out;
  assign early_reset_static_par0_go_in = wrapper_early_reset_static_par0_go_out; // @[]
  assign early_reset_static_par0_done_in = ud3_out;
  assign early_reset_static_seq_go_in = wrapper_early_reset_static_seq_go_out; // @[]
  assign early_reset_static_seq_done_in = ud4_out;
  assign early_reset_static_par1_go_in = wrapper_early_reset_static_par1_go_out; // @[]
  assign early_reset_static_par1_done_in = ud5_out;
  assign early_reset_static_seq1_go_in = wrapper_early_reset_static_seq1_go_out; // @[]
  assign early_reset_static_seq1_done_in = ud6_out;
  assign wrapper_early_reset_static_par_go_in = ~wrapper_early_reset_static_par_done_out & fsm9_out == 5'h0 &
    tdcc8_go_out; // @[]
  assign wrapper_early_reset_static_par_done_in = fsm_out == 5'h0 & signal_reg_out; // @[]
  assign wrapper_early_reset_cond00_go_in = ~wrapper_early_reset_cond00_done_out & fsm9_out == 5'h1 & tdcc8_go_out | ~
    wrapper_early_reset_cond00_done_out & fsm9_out == 5'h13 & tdcc8_go_out; // @[]
  assign wrapper_early_reset_cond00_done_in = fsm_out == 5'h0 & signal_reg_out; // @[]
  assign wrapper_early_reset_cond10_go_in = ~wrapper_early_reset_cond10_done_out & fsm9_out == 5'h3 & tdcc8_go_out | ~
    wrapper_early_reset_cond10_done_out & fsm9_out == 5'h11 & tdcc8_go_out; // @[]
  assign wrapper_early_reset_cond10_done_in = fsm_out == 5'h0 & signal_reg_out; // @[]
  assign wrapper_early_reset_static_par0_go_in = ~wrapper_early_reset_static_par0_done_out & fsm9_out == 5'h4 &
    tdcc8_go_out; // @[]
  assign wrapper_early_reset_static_par0_done_in = fsm_out == 5'h0 & signal_reg_out; // @[]
  assign wrapper_early_reset_cond20_go_in = ~wrapper_early_reset_cond20_done_out & fsm9_out == 5'h5 & tdcc8_go_out | ~
    wrapper_early_reset_cond20_done_out & fsm9_out == 5'hc & tdcc8_go_out; // @[]
  assign wrapper_early_reset_cond20_done_in = fsm_out == 5'h0 & signal_reg_out; // @[]
  assign wrapper_early_reset_static_seq_go_in = ~wrapper_early_reset_static_seq_done_out & fsm9_out == 5'h9 &
    tdcc8_go_out; // @[]
  assign wrapper_early_reset_static_seq_done_in = fsm_out == 5'h0 & signal_reg_out; // @[]
  assign wrapper_early_reset_static_par1_go_in = ~wrapper_early_reset_static_par1_done_out & fsm9_out == 5'hb &
    tdcc8_go_out; // @[]
  assign wrapper_early_reset_static_par1_done_in = fsm_out == 5'h0 & signal_reg_out; // @[]
  assign wrapper_early_reset_static_seq1_go_in = ~wrapper_early_reset_static_seq1_done_out & fsm9_out == 5'h10 &
    tdcc8_go_out; // @[]
  assign wrapper_early_reset_static_seq1_done_in = fsm_out == 5'h0 & signal_reg_out; // @[]
  assign par0_go_in = ~par0_done_out & fsm9_out == 5'h8 & tdcc8_go_out; // @[]
  assign par0_done_in = pd_out & pd0_out & pd1_out; // @[]
  assign tdcc_go_in = ~(pd_out | tdcc_done_out) & par0_go_out; // @[]
  assign tdcc_done_in = fsm0_out == 2'h2; // @[]
  assign tdcc0_go_in = ~(pd0_out | tdcc0_done_out) & par0_go_out; // @[]
  assign tdcc0_done_in = fsm1_out == 2'h2; // @[]
  assign tdcc1_go_in = ~(pd1_out | tdcc1_done_out) & par0_go_out; // @[]
  assign tdcc1_done_in = fsm2_out == 2'h2; // @[]
  assign par1_go_in = ~par1_done_out & fsm9_out == 5'ha & tdcc8_go_out; // @[]
  assign par1_done_in = pd2_out & pd3_out; // @[]
  assign tdcc2_go_in = ~(pd2_out | tdcc2_done_out) & par1_go_out; // @[]
  assign tdcc2_done_in = fsm3_out == 2'h2; // @[]
  assign tdcc3_go_in = ~(pd3_out | tdcc3_done_out) & par1_go_out; // @[]
  assign tdcc3_done_in = fsm4_out == 2'h2; // @[]
  assign par2_go_in = ~par2_done_out & fsm9_out == 5'hf & tdcc8_go_out; // @[]
  assign par2_done_in = pd4_out & pd5_out & pd6_out & pd7_out; // @[]
  assign tdcc4_go_in = ~(pd4_out | tdcc4_done_out) & par2_go_out; // @[]
  assign tdcc4_done_in = fsm5_out == 2'h2; // @[]
  assign tdcc5_go_in = ~(pd5_out | tdcc5_done_out) & par2_go_out; // @[]
  assign tdcc5_done_in = fsm6_out == 2'h2; // @[]
  assign tdcc6_go_in = ~(pd6_out | tdcc6_done_out) & par2_go_out; // @[]
  assign tdcc6_done_in = fsm7_out == 2'h2; // @[]
  assign tdcc7_go_in = ~(pd7_out | tdcc7_done_out) & par2_go_out; // @[]
  assign tdcc7_done_in = fsm8_out == 2'h2; // @[]
  assign tdcc8_go_in = go;
  assign tdcc8_done_in = fsm9_out == 5'h14; // @[]
endmodule
